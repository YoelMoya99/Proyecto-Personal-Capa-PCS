module onescount (
    general_code_group,
    rd_in,
    rd_out
    );


    // Lista de entradas y salidas
    input [9:0] general_code_group;
    input rd_in;
    output reg rd_out;

endmodule
